// This code is part of the model collection of simulatable TTL devices.
// Note this does not necessarily mean they are synthesizable!!!
//
// Copyright (C) 2022  Holger Veit (hveit01@web.de)
//
//    This program is free software; you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation; either version 3 of the License, or (at
//    your option) any later version.
//
//    This program is distributed in the hope that it will be useful, but
//    WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
//    General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, see <http://www.gnu.org/licenses/>.
//
//
// D FF with Preset/Clear
module sn74ls74(q, q_, d, clk, pre, clr);
input d, clk, pre, clr;
output q;
output q_;
reg ff;

parameter
	// TI TTL data book Vol 1, 1985
	tPLH_min=0, tPLH_typ=13, tPLH_max=25,
	tPHL_min=0, tPHL_typ=25, tPHL_max=40;

always @(clr==0)
begin
	ff <= 0;
end

always @(pre==0)
begin
	ff <= 1;
end	

always @(posedge clk)
begin
	if (clr==1 && pre==1)
		ff <= d;
end

assign #(tPLH_min:tPLH_typ:tPLH_max,
		 tPHL_min:tPHL_typ:tPHL_max)
	q  = pre==0 ? 1 : 
		 clr==0 ? 0 : ff;
assign #(tPLH_min:tPLH_typ:tPLH_max,
		 tPHL_min:tPHL_typ:tPHL_max)
	q_ = clr==0 ? 1 : 
		 pre==0 ? 0 : ~ff;

endmodule
